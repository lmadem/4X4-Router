//sequencer goal is to receive transactions from sequence and send it to driver through TLM ports

typedef uvm_sequencer #(packet) sequencer;