//crc_test_callback goal is to inject error into DUT by adding actual callback object to driver to corrupt CRC
class crc_test_callback extends uvm_test;
  //register crc_test_callback into factory
  `uvm_component_utils(crc_test_callback)
  
  virtual router_if vif;
  bit [31:0] dropped_pkt_count;
  bit [31:0] exp_pkt_count;  
  environment env;
  
  function new (string name="crc_test_callback",uvm_component parent=null);
    super.new(name, parent);
  endfunction
  
  //define extern methods
  extern virtual function void build_phase(uvm_phase phase);
  extern virtual function void end_of_elaboration_phase(uvm_phase phase);
  extern virtual task main_phase (uvm_phase phase);
  extern virtual task shutdown_phase (uvm_phase phase);
  extern virtual function void report_phase(uvm_phase phase);

endclass	
    
//Build-phase   
function void crc_test_callback::build_phase(uvm_phase phase);
  super.build_phase(phase);
  exp_pkt_count=5;
  env=environment::type_id::create("env",this);
  
  //Below shown all are environment(testbench) configurations
  //Get the physical interface from program block
  uvm_config_db#(virtual router_if)::get(this, "", "vif", vif);
  
  //set the test name for readability in the environment
  uvm_config_db#(string)::set(this, "env.*", "test_name", get_type_name());
  
  for(bit [2:0] i=1; i<=4; i++) begin
    //below are to set the physical interface to child components (drvr,iMon and oMon) 
    //Set the physical interface to Driver
    uvm_config_db#(virtual router_if.tb_mod_port)::set(this, $sformatf("env.m_agent[%0d]", i), "drvr_if", vif.tb_mod_port);
  
    //Set the physical interface to Input Monitor
    uvm_config_db#(virtual router_if.tb_mon)::set(this, $sformatf("env.m_agent[%0d]", i), "iMon_if", vif.tb_mon);
  
    //Set the physical interface to Output Monitor
    uvm_config_db#(virtual router_if.tb_mon)::set(this, $sformatf("env.s_agent[%0d]", i), "oMon_if", vif.tb_mon);
    
    //set the pkt count to be generated by sequence
    uvm_config_db#(int)::set(this, $sformatf("env.m_agent[%0d].seqr", i), "item_count", exp_pkt_count);
  end
  
  //Set the number of packets to retain in environment for the validation of test
  uvm_config_db#(int)::set(this, "env", "item_count", exp_pkt_count*4);
  
  //Below shown settings are to configure sequencer to execute particular sequence in a particular phase
  
  //configure sequencer to execute reset_sequence in reset_phase of sequencer
  uvm_config_db#(uvm_object_wrapper)::set(this, "env.m_agent[1].seqr.reset_phase", "default_sequence", reset_sequence::get_type());
  
  //configure sequencer to execute config_sequence in configure_phase of sequencer
  uvm_config_db#(uvm_object_wrapper)::set(this, "env.m_agent[1].seqr.configure_phase", "default_sequence", config_sequence::get_type());
  
  //configure sequencer to execute sa1_da1_sequence in main_phase of sequencer
  uvm_config_db#(uvm_object_wrapper)::set(this, "env.m_agent[1].seqr.main_phase", "default_sequence", crc_sequence::get_type());
  
  //configure sequencer to execute sa2_da2_sequence in main_phase of sequencer
  uvm_config_db#(uvm_object_wrapper)::set(this, "env.m_agent[2].seqr.main_phase", "default_sequence", crc_sequence::get_type());
  
  //configure sequencer to execute sa3_da3_sequence in main_phase of sequencer
  uvm_config_db#(uvm_object_wrapper)::set(this, "env.m_agent[3].seqr.main_phase", "default_sequence", crc_sequence::get_type());
  
  //configure sequencer to execute sa4_da4_sequence in main_phase of sequencer
  uvm_config_db#(uvm_object_wrapper)::set(this, "env.m_agent[4].seqr.main_phase", "default_sequence", crc_sequence::get_type());
  
  uvm_config_db#(bit)::set(this,"env","enable_report",1'b1); 

endfunction
    
//Implement end_of_elaboration_phase to add callbacks       
function void crc_test_callback::end_of_elaboration_phase(uvm_phase phase);
  //handle drv_err_cb of type err_inject_drv_cb
  crc_err_inject_drv_cb crc_drv_err_cb;
  super.end_of_elaboration_phase(phase);
  
  //Construct callback object crc_drv_err_cb
  crc_drv_err_cb = new();
  
  //Add callback object crc_drv_err_cb to driver
  uvm_callbacks #(driver, driver_callback_facade_crc)::add(this.env.m_agent[1].drvr, crc_drv_err_cb);
  
  uvm_callbacks #(driver, driver_callback_facade_crc)::add(this.env.m_agent[2].drvr, crc_drv_err_cb);
    
  uvm_callbacks #(driver, driver_callback_facade_crc)::add(this.env.m_agent[3].drvr, crc_drv_err_cb);
    
  uvm_callbacks #(driver, driver_callback_facade_crc)::add(this.env.m_agent[4].drvr, crc_drv_err_cb);

  uvm_callbacks #(driver, driver_callback_facade_crc)::display();
   
endfunction

//main phase
task crc_test_callback::main_phase(uvm_phase phase);
  uvm_objection objection;
  super.main_phase(phase);
  objection=phase.get_objection();
  objection.set_drain_time(this,2500ns);
  //The drain time is the amount of time to wait once all objections have been dropped
endtask

//Run shutdown sequence in shutdown phase to read drooped count from DUT
task crc_test_callback::shutdown_phase(uvm_phase phase);
  //Instantiate and construct shutdown sequence
  crc_shutdown_sequence seq;
  seq = crc_shutdown_sequence::type_id::create("seq", this);
  phase.raise_objection(this, "Raised objection from CRC callback test");
  //Start the shutdown seq on sequencer
  seq.start(this.env.m_agent[1].seqr);
  
  //Get the dropped count from seq which helps in deciding test pass or fail
  dropped_pkt_count = seq.dropped_pkt_count;
  phase.drop_objection(this, "Dropped objection from CRC callback test");
endtask
      
//report_phase to print test PASS or FAIL results.
function void crc_test_callback::report_phase(uvm_phase phase);
  //Check if total pkts dropped by dut equal to pkts driven into DUT 
  if(exp_pkt_count*4 != dropped_pkt_count) begin

    `uvm_info("FAIL", "****************Test FAILED******************", UVM_NONE);
    `uvm_info("FAIL","Test Failed due to packet count MIS_MATCH",UVM_NONE); 
    `uvm_info("FAIL",$sformatf("exp_pkt_count=%0d Dropped_pkt_count=%0d ",exp_pkt_count*4,dropped_pkt_count),UVM_NONE); 
    `uvm_fatal("FAIL","******************Test FAILED ************");
  end
  //Test Passed as all packets dropped by DUT.
  else begin
    `uvm_info("PASS", "******************Test PASSED ***************",UVM_NONE);
    `uvm_info("PASS",$sformatf("exp_pkt_count=%0d Dropped_pkt_count=%0d ",exp_pkt_count*4,dropped_pkt_count),UVM_NONE); 
    `uvm_info("PASS","******************************************",UVM_NONE);
  end
endfunction


