// Code your testbench here
// or browse Examples
//`include "test.sv" - This is a linear testbench, always comment it when the SV environment is ON

`include "top.sv"
`include "interface.sv"
`include "program_test.sv"




