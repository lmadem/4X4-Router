package router_pkg;
`include "header.h"
`include "packet.sv"
`include "generator.sv"
`include "driver.sv"
`include "iMonitor.sv"
`include "oMonitor.sv"
`include "scoreboard.sv"
`include "coverage.sv"
`include "generator_ext.sv"
`include "environment.sv"
endpackage
