// Code your testbench here
// or browse Examples
`include "top.sv"               //Top Module
`include "router_if.sv"         //Interface
`include "program_router_tb.sv" //Program Block 